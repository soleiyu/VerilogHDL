//lemon3 yonedu

module lemon3
(
	input	wire  [9:0]		count,  
	output wire [15:0]  	outv
);

	reg [15:0] notes [1023:0];
	assign outv = notes[count];

	initial
	begin
	notes[14] <= {8'd1, 8'd51};
	notes[15] <= {8'd1, 8'd53};
	
	notes[16] <= {8'd2, 8'd55};
	notes[17] <= {8'd1, 8'd51};
	notes[18] <= {8'd1, 8'd48};
	notes[19] <= {8'd2, 8'd0};
	notes[20] <= {8'd2, 8'd53};
	notes[21] <= {8'd2, 8'd50};
	notes[22] <= {8'd1, 8'd46};
	notes[23] <= {8'd1, 8'd43};
	notes[24] <= {8'd2, 8'd0};
	notes[25] <= {8'd2, 8'd50};
	
	notes[26] <= {8'd2, 8'd48};
	notes[27] <= {8'd1, 8'd46};
	notes[28] <= {8'd3, 8'd39};
	notes[29] <= {8'd2, 8'd46};
	notes[30] <= {8'd4, 8'd43};
	notes[31] <= {8'd2, 8'd0};
	notes[32] <= {8'd1, 8'd41};
	notes[33] <= {8'd1, 8'd43};
	
	notes[34] <= {8'd4, 8'd44};
	notes[35] <= {8'd2, 8'd51};
	notes[36] <= {8'd1, 8'd50};
	notes[37] <= {8'd1, 8'd51};
	notes[38] <= {8'd4, 8'd46};
	notes[39] <= {8'd2, 8'd44};
	notes[40] <= {8'd1, 8'd43};
	notes[41] <= {8'd1, 8'd44};
 
	notes[42] <= {8'd3, 8'd45};
	notes[43] <= {8'd1, 8'd45};
	notes[44] <= {8'd2, 8'd51};
	notes[45] <= {8'd1, 8'd50};
	notes[46] <= {8'd1, 8'd48};
	notes[47] <= {8'd4, 8'd47};
	notes[48] <= {8'd2, 8'd0};
	notes[49] <= {8'd1, 8'd51};
	notes[50] <= {8'd1, 8'd53};
	
	notes[51] <= {8'd2, 8'd55};
	notes[52] <= {8'd1, 8'd51};
	notes[53] <= {8'd1, 8'd48};
	notes[54] <= {8'd2, 8'd0};
	notes[55] <= {8'd2, 8'd53};
	notes[56] <= {8'd2, 8'd50};
	notes[57] <= {8'd1, 8'd46};
	notes[58] <= {8'd1, 8'd43};
	notes[59] <= {8'd2, 8'd0};
	notes[60] <= {8'd2, 8'd50};
	
	notes[61] <= {8'd2, 8'd48};
	notes[62] <= {8'd1, 8'd46};
	notes[63] <= {8'd3, 8'd39};
	notes[64] <= {8'd2, 8'd46};
	notes[65] <= {8'd4, 8'd43};
	notes[66] <= {8'd2, 8'd0};
	notes[67] <= {8'd1, 8'd41};
	notes[68] <= {8'd1, 8'd43};
 
	notes[69] <= {8'd4, 8'd44};
	notes[70] <= {8'd2, 8'd46};
	notes[71] <= {8'd1, 8'd44};
	notes[72] <= {8'd1, 8'd46};
	notes[73] <= {8'd2, 8'd43};
	notes[74] <= {8'd2, 8'd46};
	notes[75] <= {8'd2, 8'd51};
	notes[76] <= {8'd2, 8'd55};
	
	notes[77] <= {8'd3, 8'd53};
	notes[78] <= {8'd1, 8'd53};
	notes[79] <= {8'd3, 8'd53};
	notes[80] <= {8'd1, 8'd51};
	notes[81] <= {8'd8, 8'd51};	
	
	notes[82] <= {8'd14, 8'd0};
	notes[83] <= {8'd1, 8'd51};
	notes[84] <= {8'd1, 8'd53};
	
	notes[85] <= {8'd2, 8'd55};
	notes[86] <= {8'd1, 8'd51};
	notes[87] <= {8'd1, 8'd48};
	notes[88] <= {8'd2, 8'd0};
	notes[89] <= {8'd2, 8'd53};
	notes[90] <= {8'd2, 8'd50};
	notes[91] <= {8'd1, 8'd46};
	notes[92] <= {8'd1, 8'd43};
	notes[93] <= {8'd2, 8'd0};
	notes[94] <= {8'd2, 8'd50};
	
	notes[95] <= {8'd2, 8'd48};
	notes[96] <= {8'd1, 8'd46};
	notes[97] <= {8'd3, 8'd39};
	notes[98] <= {8'd2, 8'd46};
	notes[99] <= {8'd4, 8'd43};
	notes[100] <= {8'd2, 8'd0};
	notes[101] <= {8'd1, 8'd41};
	notes[102] <= {8'd1, 8'd43};
	
	notes[103] <= {8'd4, 8'd44};
	notes[104] <= {8'd2, 8'd51};
	notes[105] <= {8'd1, 8'd50};
	notes[106] <= {8'd1, 8'd51};
	notes[107] <= {8'd4, 8'd46};
	notes[108] <= {8'd2, 8'd44};
	notes[109] <= {8'd1, 8'd43};
	notes[110] <= {8'd1, 8'd44};
 
	notes[111] <= {8'd4, 8'd45};
	notes[112] <= {8'd2, 8'd51};
	notes[113] <= {8'd1, 8'd50};
	notes[114] <= {8'd1, 8'd48};
	notes[115] <= {8'd4, 8'd47};
	notes[116] <= {8'd2, 8'd0};
	notes[117] <= {8'd1, 8'd51};
	notes[118] <= {8'd1, 8'd53};
	
	notes[119] <= {8'd2, 8'd55};
	notes[120] <= {8'd1, 8'd51};
	notes[121] <= {8'd1, 8'd48};
	notes[122] <= {8'd2, 8'd0};
	notes[123] <= {8'd2, 8'd53};
	notes[124] <= {8'd2, 8'd50};
	notes[125] <= {8'd1, 8'd46};
	notes[126] <= {8'd1, 8'd43};
	notes[127] <= {8'd2, 8'd0};
	notes[128] <= {8'd2, 8'd50};
	
	notes[129] <= {8'd2, 8'd48};
	notes[130] <= {8'd1, 8'd46};
	notes[131] <= {8'd3, 8'd39};
	notes[132] <= {8'd2, 8'd46};
	notes[133] <= {8'd4, 8'd43};
	notes[134] <= {8'd2, 8'd0};
	notes[135] <= {8'd1, 8'd41};
	notes[136] <= {8'd1, 8'd43};
 
	notes[137] <= {8'd4, 8'd44};
	notes[138] <= {8'd2, 8'd46};
	notes[139] <= {8'd1, 8'd44};
	notes[140] <= {8'd1, 8'd46};
	notes[141] <= {8'd2, 8'd43};
	notes[142] <= {8'd2, 8'd46};
	notes[143] <= {8'd2, 8'd51};
	notes[144] <= {8'd2, 8'd55};
	
	notes[145] <= {8'd1, 8'd53};
	notes[146] <= {8'd3, 8'd53};
	notes[147] <= {8'd3, 8'd53};
	notes[148] <= {8'd1, 8'd51};
	notes[149] <= {8'd8, 8'd51};

	
	notes[150] <= {8'd3, 8'd48};
	notes[151] <= {8'd1, 8'd50};
	notes[152] <= {8'd2, 8'd51};
	notes[153] <= {8'd1, 8'd50};
	notes[154] <= {8'd1, 8'd48};
	notes[155] <= {8'd2, 8'd46};
	notes[156] <= {8'd2, 8'd55};
	notes[157] <= {8'd2, 8'd55};
	notes[158] <= {8'd2, 8'd0};
	
	notes[159] <= {8'd3, 8'd53};
	notes[160] <= {8'd1, 8'd55};
	notes[161] <= {8'd2, 8'd56};
	notes[162] <= {8'd1, 8'd55};
	notes[163] <= {8'd1, 8'd53};
	notes[164] <= {8'd2, 8'd51};
	notes[165] <= {8'd2, 8'd53};
	notes[166] <= {8'd2, 8'd46};
	notes[167] <= {8'd2, 8'd0};
	
	notes[168] <= {8'd3, 8'd44};
	notes[169] <= {8'd1, 8'd46};
	notes[170] <= {8'd2, 8'd48};
	notes[171] <= {8'd1, 8'd46};
	notes[172] <= {8'd1, 8'd44};
	notes[173] <= {8'd2, 8'd43};
	notes[174] <= {8'd2, 8'd51};
	notes[175] <= {8'd2, 8'd51};
	notes[176] <= {8'd2, 8'd51};
	
	notes[177] <= {8'd4, 8'd50};
	notes[178] <= {8'd2, 8'd48};
	notes[179] <= {8'd2, 8'd50};
	notes[180] <= {8'd4, 8'd51};
	notes[181] <= {8'd1, 8'd53};
	notes[182] <= {8'd1, 8'd55};
	notes[183] <= {8'd1, 8'd53};
	notes[184] <= {8'd1, 8'd51};
	
	
	notes[185] <= {8'd1, 8'd48};
	notes[186] <= {8'd3, 8'd51};
	notes[187] <= {8'd1, 8'd55};
	notes[188] <= {8'd3, 8'd58};
	notes[189] <= {8'd1, 8'd53};
	notes[190] <= {8'd3, 8'd51};
	notes[191] <= {8'd1, 8'd53};
	notes[192] <= {8'd1, 8'd55};
	notes[193] <= {8'd1, 8'd53};
	notes[194] <= {8'd1, 8'd51};
	
	notes[195] <= {8'd1, 8'd48};
	notes[196] <= {8'd3, 8'd51};
	notes[197] <= {8'd1, 8'd55};
	notes[198] <= {8'd3, 8'd58};
	notes[199] <= {8'd1, 8'd53};
	notes[200] <= {8'd3, 8'd51};
	notes[201] <= {8'd1, 8'd53};
	notes[202] <= {8'd1, 8'd55};
	notes[203] <= {8'd1, 8'd53};
	notes[204] <= {8'd1, 8'd51};
	
	notes[205] <= {8'd1, 8'd48};
	notes[206] <= {8'd3, 8'd51};
	notes[207] <= {8'd1, 8'd55};
	notes[208] <= {8'd2, 8'd58};
	notes[209] <= {8'd1, 8'd58};
	notes[210] <= {8'd1, 8'd60};
	notes[211] <= {8'd3, 8'd58};
	notes[212] <= {8'd1, 8'd58};
	notes[213] <= {8'd3, 8'd63};
	
	notes[214] <= {8'd1, 8'd62};
	notes[215] <= {8'd3, 8'd58};
	notes[216] <= {8'd1, 8'd55};
	notes[217] <= {8'd3, 8'd58};
	notes[218] <= {8'd4, 8'd53};
	notes[219] <= {8'd1, 8'd53};
	notes[220] <= {8'd1, 8'd55};
	notes[221] <= {8'd1, 8'd53};
	notes[222] <= {8'd1, 8'd51};
	
	notes[223] <= {8'd1, 8'd48};
	notes[224] <= {8'd3, 8'd51};
	notes[225] <= {8'd1, 8'd55};
	notes[226] <= {8'd3, 8'd58};
	notes[227] <= {8'd1, 8'd53};
	notes[228] <= {8'd2, 8'd51};
	notes[229] <= {8'd1, 8'd51};
	notes[230] <= {8'd1, 8'd51};
	notes[231] <= {8'd1, 8'd51};
	notes[232] <= {8'd1, 8'd53};
	notes[233] <= {8'd1, 8'd55};
	
	notes[234] <= {8'd1, 8'd56};
	notes[235] <= {8'd3, 8'd55};
	notes[236] <= {8'd1, 8'd53};
	notes[237] <= {8'd3, 8'd50};
	notes[238] <= {8'd4, 8'd51};
	notes[239] <= {8'd2, 8'd0};
	notes[240] <= {8'd1, 8'd51};
	notes[241] <= {8'd1, 8'd50};
	
	notes[242] <= {8'd2, 8'd48};
	notes[243] <= {8'd2, 8'd50};
	notes[244] <= {8'd2, 8'd51};
	notes[245] <= {8'd2, 8'd53};
	notes[246] <= {8'd2, 8'd51};
	notes[247] <= {8'd2, 8'd46};
	notes[248] <= {8'd1, 8'd43};
	notes[249] <= {8'd3, 8'd46};
	
	notes[250] <= {8'd1, 8'd48};
	notes[251] <= {8'd3, 8'd53};
	notes[252] <= {8'd1, 8'd50};
	notes[253] <= {8'd3, 8'd51};
	notes[254] <= {8'd4, 8'd51};
	notes[255] <= {8'd2, 8'd0};
	notes[256] <= {8'd1, 8'd51};
	notes[257] <= {8'd1, 8'd50};
	
	notes[258] <= {8'd2, 8'd48};
	notes[259] <= {8'd2, 8'd50};
	notes[260] <= {8'd2, 8'd51};
	notes[261] <= {8'd2, 8'd53};
	notes[262] <= {8'd2, 8'd51};
	notes[263] <= {8'd2, 8'd46};
	notes[264] <= {8'd1, 8'd51};
	notes[265] <= {8'd3, 8'd53};
	
	notes[266] <= {8'd1, 8'd55};
	notes[267] <= {8'd3, 8'd56};
	notes[268] <= {8'd1, 8'd53};
	notes[269] <= {8'd3, 8'd51};
	notes[270] <= {8'd6, 8'd51};

	end
	
endmodule
